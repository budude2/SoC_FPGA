`timescale 1ns / 1ps

module reaction_test_top(

    );
endmodule
