`timescale 1ns / 1ps

module state_machine
( );
endmodule
